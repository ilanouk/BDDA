�� sr Catalogi�*�<4 L listeRelationt Ljava/util/ArrayList;xpsr java.util.ArrayListx����a� I sizexp   w   sr RelationInfo��3Ǝ� I 
nbrColonneL colonnesq ~ L nomRelationt Ljava/lang/String;xp   sq ~    w   sr ColInfo���ht.�� L nomq ~ L typeq ~ xpt nomt Integerxt testsq ~    sq ~    w   sq ~ 	t nomt Integerxt testsq ~    sq ~    w   sq ~ 	t nomt Integerxt testsq ~    sq ~    w   sq ~ 	t nomt Integerxt testx