�� sr Catalogi�*�<4 L listeRelationt Ljava/util/ArrayList;xpsr java.util.ArrayListx����a� I sizexp   w   sr RelationInfow�R�ɭ� I 
nbrColonneL colonnesq ~ L headerPageIdt LPageId;L nomRelationt Ljava/lang/String;xp   sq ~    w   sr ColInfo���ht.�� L nomq ~ L typeq ~ xpt NOMt VARCHARxsr PageId��y���|L I FileIdxI PageIdxxp       t TESTx