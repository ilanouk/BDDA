�� sr Catalogi�*�<4 L listeRelationt Ljava/util/ArrayList;xpsr java.util.ArrayListx����a� I sizexp   w   sr RelationInfow�bh� I 
nbrColonneL colonnesq ~ L headerPageIdt LPageId;L nomRelationt Ljava/lang/String;xp   sq ~    w   sr ColInfo���ht.�� L nomq ~ L typeq ~ xpt nomt INTEGERxpt testsq ~    sq ~    w   sq ~ 
t nomt INTEGERxpt testsq ~    sq ~    w   sq ~ 
t nomt INTEGERxpt testsq ~    sq ~    w   sq ~ 
t nomt INTEGERx{sr  java.io.NotSerializableException(Vx �5  xr java.io.ObjectStreamExceptiond��k�9��  xr java.io.IOExceptionl�sde%�  xr java.lang.Exception��>;�  xr java.lang.Throwable��5'9w�� L causet Ljava/lang/Throwable;L detailMessaget Ljava/lang/String;[ 
stackTracet [Ljava/lang/StackTraceElement;L suppressedExceptionst Ljava/util/List;xpq ~ 	t PageIdur [Ljava.lang.StackTraceElement;F*<<�"9  xp   sr java.lang.StackTraceElementa	Ś&6݅ B formatI 
lineNumberL classLoaderNameq ~ L declaringClassq ~ L fileNameq ~ L 
methodNameq ~ L 
moduleNameq ~ L moduleVersionq ~ xp  �pt java.io.ObjectOutputStreamt ObjectOutputStream.javat writeObject0t 	java.baset 11.0.17sq ~   pq ~ q ~ t defaultWriteFieldsq ~ q ~ sq ~   �pq ~ q ~ t writeSerialDataq ~ q ~ sq ~   �pq ~ q ~ t writeOrdinaryObjectq ~ q ~ sq ~   �pq ~ q ~ q ~ q ~ q ~ sq ~   Ypq ~ q ~ t writeObjectq ~ q ~ sq ~   �pt java.util.ArrayListt ArrayList.javaq ~ q ~ q ~ sq ~ ����pt -jdk.internal.reflect.NativeMethodAccessorImplt NativeMethodAccessorImpl.javat invoke0q ~ q ~ sq ~    >pq ~ !q ~ "t invokeq ~ q ~ sq ~    +pt 1jdk.internal.reflect.DelegatingMethodAccessorImplt !DelegatingMethodAccessorImpl.javaq ~ %q ~ q ~ sq ~   6pt java.lang.reflect.Methodt Method.javaq ~ %q ~ q ~ sq ~   �pt java.io.ObjectStreamClasst ObjectStreamClass.javat invokeWriteObjectq ~ q ~ sq ~   �pq ~ q ~ q ~ q ~ q ~ sq ~   �pq ~ q ~ q ~ q ~ q ~ sq ~   �pq ~ q ~ q ~ q ~ q ~ sq ~   pq ~ q ~ q ~ q ~ q ~ sq ~   �pq ~ q ~ q ~ q ~ q ~ sq ~   �pq ~ q ~ q ~ q ~ q ~ sq ~   �pq ~ q ~ q ~ q ~ q ~ sq ~   Ypq ~ q ~ q ~ q ~ q ~ sq ~    .t appt Catalogt Catalog.javat saveppsq ~    q ~ 9q ~ :q ~ ;t Finishppsq ~    	q ~ 9t TestCatalogt TestCatalog.javat addRelationTestppsq ~    q ~ 9q ~ @q ~ At mainppsr java.util.Collections$EmptyListz��<���  xpx